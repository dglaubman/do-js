10% share of unlimited xs 0