100% share of 1000000 xs 1000000