100% share of 10000 xs 10000