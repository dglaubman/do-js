50% share of 20000 xs 5000