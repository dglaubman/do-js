100% share of 10000000 xs 20000000