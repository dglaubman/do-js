100% share of 1000 xs 1000