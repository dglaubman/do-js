100% share of unlimited xs 1000