50% share of 50000000 xs 0