100% share of 20000000 xs 15000000