100% share of 20000000 xs 5000000