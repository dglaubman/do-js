20% share of 5000 xs 1000