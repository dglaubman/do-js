90% share of unlimited xs 500