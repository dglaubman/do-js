100% share of 4000000 xs 1000000